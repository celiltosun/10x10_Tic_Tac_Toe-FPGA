////////////////////////////////////////////////////////////////////////////////////////////////////////
// Middle East Technical University Electrical and Electronical Engineering 2022-2023 Junior Year Endterm Project
// FPGA Implementation of 2D Turn Based Strategy Game(10x10 Scaled Tic Tac Toe) on VGA Display
// Created by: Ahmet Alperen Tekin & Ali Bora Metin & Arman Özcan & Celil Tosun
///////////////////////////////////////////////////////////////////////////////////////////////////////

//-----------------VGA Display Part---------------------------------
module vga_display(divided_clk, V_Sync, H_Sync, board, R_out, G_out, B_out, turn, wld, roundcount, triwincount, circwincount, error);

	input wire divided_clk;
	input wire [299:0] board;
	input wire [4:0] roundcount;
	output reg V_Sync;
	output reg H_Sync; 
	output reg [7:0] R_out;
	output reg [7:0] G_out;
	output reg [7:0] B_out;
	input wire turn;
	input wire [1:0] wld;
	input wire [3:0] triwincount;
	input wire [3:0] circwincount;
	input wire error;
	
	reg [6335:0] triangle_won;
	reg [6335:0] draw;
	reg [19007:0] circles_turn_symbol;
	reg [19007:0] trig_turn_symbol;
	reg [6335:0] circles_won;
	reg [468:0] total_moves;
	reg [188:0] wins;
	reg [223:0] error_msg;
	reg [34:0] zero;
	reg [34:0] one;
	reg [34:0] two;
	reg [34:0] three;
	reg [34:0] four;
	reg [34:0] five;
	reg [34:0] six;
	reg [34:0] seven;
	reg [34:0] eight;
	reg [34:0] nine;
	
	
	reg [9:0] V_count;
	reg [9:0] H_count;
	
	reg in_display;
	reg in_grid_borders;
	reg counts_in_cell_range;
	wire [4:0] i;
	wire [4:0] j;
	
	parameter H_SYNC = 95; // 95
	parameter H_FRONT = 47; // 47
	parameter H_DISP = 635; // 635
	parameter H_BACK = 15; // 15
	
	parameter V_SYNC = 2; // 2
	parameter V_FRONT = 10; // 10
	parameter V_DISP = 480; // 480
	parameter V_BACK = 33; // 33
	
	parameter LIN_THCK = 2; // Grid Line Thickness
	parameter H_CELL_THCK = (H_DISP - 11*LIN_THCK - 2*H_SPAC)/10;
	parameter V_CELL_THCK = (V_DISP - 11*LIN_THCK - V_TOP_SPAC - V_BOT_SPAC)/10;
	parameter V_TOP_SPAC = 100;
	parameter V_BOT_SPAC = 50;
	parameter H_SPAC = 100;
	
	wire [7:0] R_circ;
	wire [7:0] G_circ;
	wire [7:0] B_circ;
	
	wire [7:0] R_trig;
	wire [7:0] G_trig;
	wire [7:0] B_trig;
	
	initial begin
		V_count <= 10'b0000000000; // counts up to 525
		H_count <= 10'b0000000000; // counts up to 792 
		//Texts on display with 6336 bits
		triangle_won <= 6336'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000011000011001111000000101111000111000111100000000100000100010011100000010001110000101000000000000100001000100111000101000000000101010111100011100001000000000011100011100100000100010111100011100000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000011000011001000100000101000101000101000100000000111100100010001000011110000100001010100000000000100001000101000101010100000000101010100010000010001000000000000010001000111100100010100010001000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000101111001000101000100000000100010100010001000100010000100001010100000000000000001000101000101010100000000101010111100111110001000000000111110001000100010100010111100001000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100101001101000001000101001100000000100010100110001000100010000100001010100000000000100001001101000101010100000000101010100000100010001000000000100010001000100010100110100000001000100110001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000110100111000111000110100000000011100011010001100011110000110001000100000000000100000110100111001000100000000010110011100011100001000000000011100001000011100011010011100001100011010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000001000100000000000100000000000000001000100000000000000000000000000001000000000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000001000000000000100001000100000000000100000000000000001000100000000000000000000000000111110000000000000001100000000000000000000001000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		draw <= 6336'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101111000000101111000111000111100010000010001011100000101110010100001000101001111000001000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000101000101000101000100011110010001001000111100100101010001001010101001000001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000101111001000101000100010001010001001001000100100101010000001010101111000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100101001101000001000101001100010001010011001001000100100101010001001000101000010011010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000110100111000000000110100001110001101001100111100110100010001001000100111001101010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000111000000100000000000000000000000000000100010001000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000001000000000100100010001000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		circles_turn_symbol <= 19008'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000011000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000110000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000001100000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000011000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000110000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000001100000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000011000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000110000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000001100000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000011000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000110000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000001100000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000011111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		trig_turn_symbol <= 19008'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000110000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000001100000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000010000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010000000000000000011111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000110000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000001100000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000011000000000000000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000010000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000001111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; 
		circles_won <= 6336'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000011000011001111000000101111000111000111100000000100000100010011100000010001110000101000000000000100001000100111000101000000000101010111100011100001000000000011110011100011100011100000010011100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000011000011001000100000101000101000101000100000000111100100010001000011110000100001010100000000000100001000101000101010100000000101010100010000010001000000000100000000010001000100010000010001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000101111001000101000100000000100010100010001000100010000100001010100000000000000001000101000101010100000000101010111100111110001000000000011100111110001000000010000010001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100101001101000001000101001100000000100010100110001000100010000100001010100000000000100001001101000101010100000000101010100000100010001000000000000010100010001000000010100110001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000110100111000111000110100000000011100011010001100011110000110001000100000000000100000110100111001000100000000010110011100011100001000000000011100011100001000011100011010001100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000001000100000000000100000000000000001000100000000000000000000000000001000000000000000000000001000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000001000000000000100001000100000000000100000000000000001000100000000000000000000000000111110000000000000000000001100000000000000001000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		total_moves <= 469'b0000011110011100001000011100101010000001110011110001100001110000100110010000000001001010010001010101000000010001000101001001000100010011000111001111101000101000101010100000001000111100000100100010001000000000010100010100010100010101010000000100010000000010010001000100110001110001110010001001110001011000000010000111000011100111000010011000000000000000000000000000000000000001000000000000100000000001000000000000000000000000000000000000000000110000000000010000000011111;
		wins <= 189'b000001111010001001110001010110010000010001000100010101110001110010001000100010101000000001010011000100010101110001110001101000110010001110000000000000000000010001000000000000000000100010001;
		error_msg <= 224'b10000001001110000001000001011111100000010100010000010000010000010000000101000100000100000100000110010011010001010011010011001111100011010011100011010011010000011000000000000000000000000000000110000000000000000000000000011111;
		zero <= 35'b01110100011001110101110011000101110;
		one <= 35'b01110001000010000100001000011000100;
		two <= 35'b11111000100010001000100001000101110;
		three <= 35'b01110100011000001000001000100011111;
		four <= 35'b01000010001111101001010100110001000;
		five <= 35'b01110100011000010000011110000111111;
		six <= 35'b01110100011000101111000010001001100;
		seven <= 35'b00010000100001000100010001000011111;
		eight <= 35'b01110100011000101110100011000101110;
		nine <= 35'b00110010001000011110100011000101110;
		
	
	end
	
	count_to_index cti (.H_count(H_count), .V_count(V_count), .i(i), .j(j));
	
	draw_circle(.H_count(H_count), .V_count(V_count), .i(i), .j(j), .R_out(R_circ), .G_out(G_circ), .B_out(B_circ));
	draw_trig(.H_count(H_count), .V_count(V_count), .i(i), .j(j), .R_out(R_trig), .G_out(G_trig), .B_out(B_trig));
	always @(posedge divided_clk) begin
		// horizontal & vertical sync counters that count at every positive clock edge
		if(H_count < H_SYNC + H_FRONT + H_DISP + H_BACK) begin // 792
			H_count <= H_count + 1;
		end
		
		else begin
			H_count <= 10'b0000000000;
			if(V_count < V_SYNC + V_FRONT + V_DISP + V_BACK) begin // 525
				V_count <= V_count + 1;
			end
			
			else begin
				V_count <= 10'b0000000000;
			end
		end
		
		// timing counters are set. Now, output signals are toggled according to the counters
		H_Sync <= (H_count >  0 && H_count <= H_SYNC) ? 0 : 1;
		V_Sync <= (V_count >  0 && V_count <= V_SYNC) ?  0 : 1;
		
		in_display = (H_count > H_SYNC + H_FRONT && H_count <=H_SYNC + H_FRONT + H_DISP &&
			V_count > V_SYNC + V_FRONT && V_count <= V_SYNC + V_FRONT + V_DISP);
		
		in_grid_borders = (V_count > V_SYNC + V_FRONT + V_TOP_SPAC &&
				V_count < V_SYNC + V_FRONT + LIN_THCK + V_TOP_SPAC && 
				H_count > H_SYNC + H_FRONT + H_SPAC &&
				H_count < H_SYNC + H_FRONT + H_DISP - H_SPAC) // TOP GRID BORDER
				
				||(H_count > H_SYNC + H_FRONT + H_SPAC && H_count < H_SYNC + H_FRONT + LIN_THCK + H_SPAC &&
				V_count > V_SYNC + V_FRONT + V_TOP_SPAC && 
				V_count < V_SYNC + V_FRONT + V_DISP - V_BOT_SPAC) || // LEFT GRID BORDER
				
				((H_count > H_SYNC + H_FRONT + H_SPAC + 1*LIN_THCK + 1*H_CELL_THCK && H_count <= H_SYNC + H_FRONT + 
				2*LIN_THCK + 1*H_CELL_THCK + H_SPAC) ||// periodic horizontal grid borders
				(V_count > V_SYNC + V_FRONT + 1*LIN_THCK + 1*V_CELL_THCK + V_TOP_SPAC&& 
				V_count < V_SYNC + V_FRONT + 2*LIN_THCK + 1*V_CELL_THCK + V_TOP_SPAC)  || 
				
				(H_count > H_SYNC + H_FRONT + H_SPAC + 2*LIN_THCK + 2*H_CELL_THCK && H_count <= H_SYNC + H_FRONT + 
				3*LIN_THCK + 2*H_CELL_THCK + H_SPAC) ||// periodic horizontal grid borders
				(V_count > V_SYNC + V_FRONT + 2*LIN_THCK + 2*V_CELL_THCK + V_TOP_SPAC&& 
				V_count < V_SYNC + V_FRONT + 3*LIN_THCK + 2*V_CELL_THCK + V_TOP_SPAC)  || 
				
				(H_count > H_SYNC + H_FRONT + H_SPAC + 3*LIN_THCK + 3*H_CELL_THCK && H_count <= H_SYNC + H_FRONT + 
				4*LIN_THCK + 3*H_CELL_THCK + H_SPAC) ||// periodic horizontal grid borders
				(V_count > V_SYNC + V_FRONT + 3*LIN_THCK + 3*V_CELL_THCK + V_TOP_SPAC&& 
				V_count < V_SYNC + V_FRONT + 4*LIN_THCK + 3*V_CELL_THCK + V_TOP_SPAC)  || 
				
				(H_count > H_SYNC + H_FRONT + H_SPAC + 4*LIN_THCK + 4*H_CELL_THCK && H_count <= H_SYNC + H_FRONT + 
				5*LIN_THCK + 4*H_CELL_THCK + H_SPAC) ||// periodic horizontal grid borders
				(V_count > V_SYNC + V_FRONT + 4*LIN_THCK + 4*V_CELL_THCK + V_TOP_SPAC&& 
				V_count < V_SYNC + V_FRONT + 5*LIN_THCK + 4*V_CELL_THCK + V_TOP_SPAC)  || 
				
				(H_count > H_SYNC + H_FRONT + H_SPAC + 5*LIN_THCK + 5*H_CELL_THCK && H_count <= H_SYNC + H_FRONT + 
				6*LIN_THCK + 5*H_CELL_THCK + H_SPAC) ||// periodic horizontal grid borders
				(V_count > V_SYNC + V_FRONT + 5*LIN_THCK + 5*V_CELL_THCK + V_TOP_SPAC&& 
				V_count < V_SYNC + V_FRONT + 6*LIN_THCK + 5*V_CELL_THCK + V_TOP_SPAC)  || 
				
				(H_count > H_SYNC + H_FRONT + H_SPAC + 6*LIN_THCK + 6*H_CELL_THCK && H_count <= H_SYNC + H_FRONT + 
				7*LIN_THCK + 6*H_CELL_THCK + H_SPAC) ||// periodic horizontal grid borders
				(V_count > V_SYNC + V_FRONT + 6*LIN_THCK + 6*V_CELL_THCK + V_TOP_SPAC&& 
				V_count < V_SYNC + V_FRONT + 7*LIN_THCK + 6*V_CELL_THCK + V_TOP_SPAC)  || 
				
				(H_count > H_SYNC + H_FRONT + H_SPAC + 7*LIN_THCK + 7*H_CELL_THCK && H_count <= H_SYNC + H_FRONT + 
				8*LIN_THCK + 7*H_CELL_THCK + H_SPAC) ||// periodic horizontal grid borders
				(V_count > V_SYNC + V_FRONT + 7*LIN_THCK + 7*V_CELL_THCK + V_TOP_SPAC&& 
				V_count < V_SYNC + V_FRONT + 8*LIN_THCK + 7*V_CELL_THCK + V_TOP_SPAC)  || 
				
				(H_count > H_SYNC + H_FRONT + H_SPAC + 8*LIN_THCK + 8*H_CELL_THCK && H_count <= H_SYNC + H_FRONT + 
				9*LIN_THCK + 8*H_CELL_THCK + H_SPAC) ||// periodic horizontal grid borders
				(V_count > V_SYNC + V_FRONT + 8*LIN_THCK + 8*V_CELL_THCK + V_TOP_SPAC&& 
				V_count < V_SYNC + V_FRONT + 9*LIN_THCK + 8*V_CELL_THCK + V_TOP_SPAC)  || 
				
				(H_count > H_SYNC + H_FRONT + H_SPAC + 9*LIN_THCK + 9*H_CELL_THCK && H_count <= H_SYNC + H_FRONT + 
				10*LIN_THCK + 9*H_CELL_THCK + H_SPAC) ||// periodic horizontal grid borders
				(V_count > V_SYNC + V_FRONT + 9*LIN_THCK + 9*V_CELL_THCK + V_TOP_SPAC&& 
				V_count < V_SYNC + V_FRONT + 10*LIN_THCK + 9*V_CELL_THCK + V_TOP_SPAC)  ||
				
				(H_count > H_SYNC + H_FRONT + H_SPAC + 10*LIN_THCK + 10*H_CELL_THCK && H_count <= H_SYNC + H_FRONT + 
				11*LIN_THCK + 10*H_CELL_THCK + H_SPAC) ||// periodic horizontal grid borders
				(V_count > V_SYNC + V_FRONT + 10*LIN_THCK + 10*V_CELL_THCK + V_TOP_SPAC&& 
				V_count < V_SYNC + V_FRONT + 11*LIN_THCK + 10*V_CELL_THCK + V_TOP_SPAC))
			
				&& (V_count > V_SYNC + V_FRONT + V_TOP_SPAC + LIN_THCK && 
						V_count < V_SYNC + V_FRONT + V_DISP - V_BOT_SPAC && 
						
						H_count > H_SYNC + H_FRONT + H_SPAC + LIN_THCK &&
						H_count < H_SYNC + H_FRONT + H_DISP - H_SPAC)? 1 : 0;			
				
		
		if(in_display && ~in_grid_borders) begin			
			if (~(i == 0 || j == 0))begin
				case (board[30*(i-1) + 3*(j-1)+: 3])					
					
					3'b010 : begin
						R_out <= R_circ;//Red_square;
						G_out <= G_circ;//Green_square;
						B_out <= B_circ;//Blue_square;

					end
					
					3'b000 : begin
						R_out <= 8'b00000000;
						G_out <= 8'b00000000;
						B_out <= 8'b00000000;
					end
					
					
					3'b110 : begin
						R_out <= 8'b11111111;
						G_out <= 8'b00000000;
						B_out <= 8'b00000000;
					end
					
					3'b100 : begin
						R_out <= R_trig;
						G_out <= G_trig;
						B_out <= B_trig;
					end
					
					default : begin
						R_out <= 8'b10000110;
						G_out <= 8'b10000000;
						B_out <= 8'b10011000;
					end
				endcase
			end
			
			else if(V_count > V_SYNC + V_FRONT + 35 && V_count <= V_SYNC + V_FRONT + 43) begin
				case(wld)
					2'b01 : begin
						R_out <= triangle_won[(V_count - V_SYNC - V_FRONT - 36)*792 + H_count] ? 8'b11111111 : 8'b00000000;
						G_out <= triangle_won[(V_count - V_SYNC - V_FRONT - 36)*792 + H_count] ? 8'b11111111 : 8'b00000000;
						B_out <= triangle_won[(V_count - V_SYNC - V_FRONT - 36)*792 + H_count] ? 8'b11111111 : 8'b00000000;

					end
				
					2'b10 : begin
						R_out <= circles_won[(V_count - V_SYNC - V_FRONT - 36)*792 + H_count] ? 8'b11111111 : 8'b00000000;
						G_out <= circles_won[(V_count - V_SYNC - V_FRONT - 36)*792 + H_count] ? 8'b11111111 : 8'b00000000;
						B_out <= circles_won[(V_count - V_SYNC - V_FRONT - 36)*792 + H_count] ? 8'b11111111 : 8'b00000000;
					end
				
					2'b11 : begin
						R_out <= draw[(V_count - V_SYNC - V_FRONT - 36)*792 + H_count] ? 8'b11111111 : 8'b00000000;
						G_out <= draw[(V_count - V_SYNC - V_FRONT - 36)*792 + H_count] ? 8'b11111111 : 8'b00000000;
						B_out <= draw[(V_count - V_SYNC - V_FRONT - 36)*792 + H_count] ? 8'b11111111 : 8'b00000000;
					end
				
					default : begin
						R_out <= 8'b00000000;
						G_out <= 8'b00000000;
						B_out <= 8'b00000000;
					end	
				endcase
			end
		
			else if(V_count > V_SYNC + V_FRONT + 63 && V_count <= V_SYNC + V_FRONT + 87) begin
				case(turn)
					1'b0 : begin
						R_out <= trig_turn_symbol[(V_count - V_SYNC - V_FRONT - 64)*792 + H_count] ? 8'b11111111 : 8'b00000000;
						G_out <= trig_turn_symbol[(V_count - V_SYNC - V_FRONT - 64)*792 + H_count] ? 8'b11111111 : 8'b00000000;
						B_out <= trig_turn_symbol[(V_count - V_SYNC - V_FRONT - 64)*792 + H_count] ? 8'b11111111 : 8'b00000000;
					end
			
					1'b1 : begin
						R_out <= circles_turn_symbol[(V_count - V_SYNC - V_FRONT - 64)*792 + H_count] ? 8'b11111111 : 8'b00000000;
						G_out <= circles_turn_symbol[(V_count - V_SYNC - V_FRONT - 64)*792 + H_count] ? 8'b11111111 : 8'b00000000;
						B_out <= circles_turn_symbol[(V_count - V_SYNC - V_FRONT - 64)*792 + H_count] ? 8'b11111111 : 8'b00000000;
					end
					
					default : begin
						R_out <= circles_turn_symbol[(V_count - V_SYNC - V_FRONT - 64)*792 + H_count] ? 8'b11111111 : 8'b00000000;
						G_out <= circles_turn_symbol[(V_count - V_SYNC - V_FRONT - 64)*792 + H_count] ? 8'b11111111 : 8'b00000000;
						B_out <= circles_turn_symbol[(V_count - V_SYNC - V_FRONT - 64)*792 + H_count] ? 8'b11111111 : 8'b00000000;
					end
				endcase
			end			
			
			// total moves
			else if(V_count > V_SYNC + V_FRONT + V_TOP_SPAC + 11*LIN_THCK + 10*V_CELL_THCK + 15 && 
			V_count <= V_SYNC + V_FRONT + V_TOP_SPAC + 11*LIN_THCK + 10*V_CELL_THCK + 22 && 
			H_count > H_SYNC + H_FRONT + 50 && H_count <= H_SYNC + H_FRONT + 50 + 67) begin
				
				R_out <= total_moves[H_count - H_SYNC - H_FRONT - 51 + 67*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
				G_out <= total_moves[H_count - H_SYNC - H_FRONT - 51 + 67*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
				B_out <= total_moves[H_count - H_SYNC - H_FRONT - 51 + 67*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
			end
			
			// total move MSD
			else if(V_count > V_SYNC + V_FRONT + V_TOP_SPAC + 11*LIN_THCK + 10*V_CELL_THCK + 15 && 
			V_count <= V_SYNC + V_FRONT + V_TOP_SPAC + 11*LIN_THCK + 10*V_CELL_THCK + 22 && 
			H_count > H_SYNC + H_FRONT + 50 + 70 && H_count <= H_SYNC + H_FRONT + 50 + 70 + 5) begin
				
				if(roundcount < 10) begin
					R_out <= zero[H_count - H_SYNC - H_FRONT - 50 - 71 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					G_out <= zero[H_count - H_SYNC - H_FRONT - 50 - 71 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					B_out <= zero[H_count - H_SYNC - H_FRONT - 50 - 71 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;

				end
				
				else if (roundcount >= 10 && roundcount < 20) begin
					R_out <= one[H_count - H_SYNC - H_FRONT - 50 - 71 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					G_out <= one[H_count - H_SYNC - H_FRONT - 50 - 71 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					B_out <= one[H_count - H_SYNC - H_FRONT - 50 - 71 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;

				end
				
				else begin
					R_out <= two[H_count - H_SYNC - H_FRONT - 50 - 71 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					G_out <= two[H_count - H_SYNC - H_FRONT - 50 - 71 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					B_out <= two[H_count - H_SYNC - H_FRONT - 50 - 71 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;

				end
				
			end

			
			//total move LSD
			else if (V_count > V_SYNC + V_FRONT + V_TOP_SPAC + 11*LIN_THCK + 10*V_CELL_THCK + 15 && 
			V_count <= V_SYNC + V_FRONT + V_TOP_SPAC + 11*LIN_THCK + 10*V_CELL_THCK + 22 &&
			H_count > H_SYNC + H_FRONT + 50 + 70 + 10 && H_count <= H_SYNC + H_FRONT + 50 + 70 + 15) begin
				
				if(roundcount == 0 || roundcount - 10 == 0 || roundcount - 20 == 0) begin
					R_out <= zero[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					G_out <= zero[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					B_out <= zero[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
				end
				else if(roundcount == 1 || roundcount - 10 == 1 || roundcount - 20 == 1) begin
					R_out <= one[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					G_out <= one[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					B_out <= one[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
				end
				else if(roundcount == 2 || roundcount - 10 == 2 || roundcount - 20 == 2) begin
					R_out <= two[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					G_out <= two[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					B_out <= two[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
				end
				else if(roundcount == 3 || roundcount - 10 == 3 || roundcount - 20 == 3) begin
					R_out <= three[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					G_out <= three[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					B_out <= three[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
				end
				else if(roundcount == 4 || roundcount - 10 == 4 || roundcount - 20 == 4) begin
					R_out <= four[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					G_out <= four[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					B_out <= four[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
				end
				else if(roundcount == 5 || roundcount - 10 == 5 || roundcount - 20 == 5) begin
					R_out <= five[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					G_out <= five[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					B_out <= five[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
				end
				else if(roundcount == 6 || roundcount - 10 == 6) begin
					R_out <= six[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					G_out <= six[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					B_out <= six[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
				end
				else if(roundcount == 7 || roundcount - 10 == 7) begin
					R_out <= seven[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					G_out <= seven[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					B_out <= seven[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
				end
				else if(roundcount == 8 || roundcount - 10 == 8) begin
					R_out <= eight[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					G_out <= eight[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					B_out <= eight[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
				end
				else begin
					R_out <= nine[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					G_out <= nine[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
					B_out <= nine[H_count - H_SYNC - H_FRONT - 50 - 81 + 5*(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - 11*LIN_THCK - 10*V_CELL_THCK - 16)] ? 8'b11111111 : 8'b00000000;
				end
			end
			
			// error message
			else if(V_count > V_SYNC + V_FRONT + 44 && V_count <= V_SYNC + V_FRONT + 51 && 
			H_count > 300 && H_count <= 332) begin
				R_out <= (error && error_msg[32*(V_count - V_SYNC - V_FRONT - 45) + H_count - 301]) ? 8'b11111111: 8'b00000000;
				G_out <= (error && error_msg[32*(V_count - V_SYNC - V_FRONT - 45) + H_count - 301]) ? 8'b11111111: 8'b00000000;
				B_out <= (error && error_msg[32*(V_count - V_SYNC - V_FRONT - 45) + H_count - 301]) ? 8'b11111111: 8'b00000000;
			end
			//wins
			else if(V_count > V_SYNC + V_FRONT + 55 && V_count <= V_SYNC + V_FRONT + 62 &&
			H_count > 550 && H_count <= 550 + 27) begin
				
				R_out <= wins[H_count - 551 + 27*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
				G_out <= wins[H_count - 551 + 27*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
				B_out <= wins[H_count - 551 + 27*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
			end
			
			// win counts for triangle
			else if(V_count > V_SYNC + V_FRONT + 55 && V_count <= V_SYNC + V_FRONT + 62 &&
			H_count > 550 + 27 + 20 && H_count <= 550 + 27 + 20 + 5) begin
				if(triwincount == 0) begin
					R_out <= zero[H_count - 550 - 27 - 21 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
					G_out <= zero[H_count - 550 - 27 - 21 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
					B_out <= zero[H_count - 550 - 27 - 21 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
				end
				else if(triwincount == 1) begin
					R_out <= one[H_count - 550 - 27 - 21 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
					G_out <= one[H_count - 550 - 27 - 21 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
					B_out <= one[H_count - 550 - 27 - 21 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
				end
				else if(triwincount == 2) begin
					R_out <= two[H_count - 550 - 27 - 21 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
					G_out <= two[H_count - 550 - 27 - 21 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
					B_out <= two[H_count - 550 - 27 - 21 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
				end
				else if(triwincount == 3) begin
					R_out <= three[H_count - 550 - 27 - 21 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
					G_out <= three[H_count - 550 - 27 - 21 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
					B_out <= three[H_count - 550 - 27 - 21 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
				end
			end

			// win counts for circle
			else if(V_count > V_SYNC + V_FRONT + 55 && V_count <= V_SYNC + V_FRONT + 62 &&
			H_count > 550 + 27 + 55 && H_count <= 550 + 27 + 55 + 5) begin
				if(circwincount == 0) begin
					R_out <= zero[H_count - 550 - 27 - 56 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
					G_out <= zero[H_count - 550 - 27 - 56 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
					B_out <= zero[H_count - 550 - 27 - 56 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
				end
				else if(circwincount == 1) begin
					R_out <= one[H_count - 550 - 27 - 56 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
					G_out <= one[H_count - 550 - 27 - 56 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
					B_out <= one[H_count - 550 - 27 - 56 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
				end
				else if(circwincount == 2) begin
					R_out <= two[H_count - 550 - 27 - 56 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
					G_out <= two[H_count - 550 - 27 - 56 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
					B_out <= two[H_count - 550 - 27 - 56 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
				end
				else if(circwincount == 3) begin
					R_out <= three[H_count - 550 - 27 - 56 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
					G_out <= three[H_count - 550 - 27 - 56 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
					B_out <= three[H_count - 550 - 27 - 56 + 5*(V_count - V_SYNC - V_FRONT - 56)] ? 8'b11111111 : 8'b00000000;
				end
			end

			else begin
				R_out <= 8'b00000000;
				G_out <= 8'b00000000;
				B_out <= 8'b00000000;
			end
		end
		
		else if(in_display && in_grid_borders) begin
			R_out <= 8'b11111111;
			G_out <= 8'b11111111;
			B_out <= 8'b11111111;
		end
		

		else begin
			R_out<= 8'b00000000;
			G_out<= 8'b00000000;
			B_out<= 8'b00000000;
		end
	
	end
	
endmodule

// -------------------------------------Clock Dividing to 25Mhz from 50 Mhz--------------------------------------------------------------------
module clock_divider(clk, divided_clk);

	input wire clk;
	output reg divided_clk;

	initial begin
		divided_clk = 0;
	end

	always @(posedge clk) begin
		divided_clk = ~divided_clk;
	end

endmodule

// -----------------------------10x10 Square Drawing-------------------------------------------------------------------------
module count_to_index(H_count, V_count, i, j);
	input wire [9:0] H_count;
	input wire [9:0] V_count;
	output reg [4:0] i;
	output reg [4:0] j;
	
	parameter H_SYNC = 95; // 95
	parameter H_FRONT = 47; // 47
	parameter H_DISP = 635; // 635
	parameter H_BACK = 15; // 15
	
	parameter V_SYNC = 2; // 2
	parameter V_FRONT = 10; // 10
	parameter V_DISP = 480; // 480
	parameter V_BACK = 33; // 33
	
	parameter LIN_THCK = 2; // Grid Line Thickness
	parameter H_CELL_THCK = (H_DISP - 11*LIN_THCK - 2*H_SPAC)/10;
	parameter V_CELL_THCK = (V_DISP - 11*LIN_THCK - V_TOP_SPAC - V_BOT_SPAC)/10;
	parameter V_TOP_SPAC = 100;
	parameter V_BOT_SPAC = 50;
	parameter H_SPAC = 100;
	
	integer k;
	
	always @ (*) begin
		i = 0;
		j = 0;
		for(k = 1; k < 11; k = k + 1) begin
		
			i = (H_count > H_SYNC + H_FRONT + H_SPAC + k*LIN_THCK + (k-1)* H_CELL_THCK && 
			H_count < H_SYNC + H_FRONT + H_SPAC + k*LIN_THCK + k*H_CELL_THCK) ? k : i;
			
		
			j = (V_count > V_SYNC + V_FRONT + V_TOP_SPAC + k*LIN_THCK + (k - 1)* V_CELL_THCK && 
			V_count < V_SYNC + V_FRONT + V_TOP_SPAC + k*V_CELL_THCK + k*LIN_THCK) ? k : j;
		end		
	end
	
endmodule

//--------------------------Triangle Drawing-----------------------------------------------------

module draw_trig(H_count, V_count, i, j, R_out, G_out, B_out);
	input wire [9:0] H_count;
	input wire [9:0] V_count;
	input wire [4:0] i;
	input wire [4:0] j;
	
	output reg [7:0] R_out;
	output reg [7:0] G_out;
	output reg [7:0] B_out;
	
	parameter H_SYNC = 95; // 95
	parameter H_FRONT = 47; // 47
	parameter H_DISP = 635; // 635
	parameter H_BACK = 15; // 15
	
	parameter V_SYNC = 2; // 2
	parameter V_FRONT = 10; // 10
	parameter V_DISP = 480; // 480
	parameter V_BACK = 33; // 33
	
	parameter LIN_THCK = 2; // Grid Line Thickness
	parameter H_CELL_THCK = (H_DISP - 11*LIN_THCK - 2*H_SPAC)/10;
	parameter V_CELL_THCK = (V_DISP - 11*LIN_THCK - V_TOP_SPAC - V_BOT_SPAC)/10;
	parameter V_TOP_SPAC = 100;
	parameter V_BOT_SPAC = 50;
	parameter H_SPAC = 100;
	
	reg in_cell;
	reg write_trig;
	always @(posedge H_count) begin
		
		in_cell = (H_count > H_SYNC + H_FRONT + H_SPAC + i*LIN_THCK + (i-1)* H_CELL_THCK &&
			H_count < H_SYNC + H_FRONT + H_SPAC + i*(LIN_THCK + H_CELL_THCK) &&
			V_count > V_SYNC + V_FRONT + V_TOP_SPAC + j*LIN_THCK + (j-1)* V_CELL_THCK &&
			V_count < V_SYNC + V_FRONT + V_TOP_SPAC + j*(LIN_THCK + V_CELL_THCK)) ? 1 : 0;
		
		write_trig = (in_cell &&
			H_count - H_SYNC - H_FRONT - H_SPAC - i*LIN_THCK - (i-1)*H_CELL_THCK <
			V_count - V_SYNC - V_FRONT - V_TOP_SPAC - j*LIN_THCK - (j-1)*V_CELL_THCK) ? 1 : 0;
		
		R_out <= write_trig ? 8'b00000000 : 8'b00000000;
		G_out <= write_trig ? 8'b11111111 : 8'b00000000;
		B_out <= write_trig ? 8'b00000000 : 8'b00000000;
		
	end
	
endmodule

// ----------------------------Circle Drawing--------------------------------------------------

module draw_circle(H_count, V_count, i, j, R_out, G_out, B_out);
	input wire [9:0] H_count;
	input wire [9:0] V_count;
	input wire [4:0] i;
	input wire [4:0] j;
	
	output reg [7:0] R_out;
	output reg [7:0] G_out;
	output reg [7:0] B_out;
	
	parameter H_SYNC = 95; // 95
	parameter H_FRONT = 47; // 47
	parameter H_DISP = 635; // 635
	parameter H_BACK = 15; // 15
	
	parameter V_SYNC = 2; // 2
	parameter V_FRONT = 10; // 10
	parameter V_DISP = 480; // 480
	parameter V_BACK = 33; // 33
	
	parameter LIN_THCK = 2; // Grid Line Thickness
	parameter H_CELL_THCK = (H_DISP - 11*LIN_THCK - 2*H_SPAC)/10;
	parameter V_CELL_THCK = (V_DISP - 11*LIN_THCK - V_TOP_SPAC - V_BOT_SPAC)/10;
	parameter V_TOP_SPAC = 100;
	parameter V_BOT_SPAC = 50;
	parameter H_SPAC = 100;
	

	
	reg [9:0] H_dist;
	reg [9:0] V_dist;
	reg in_cell;
	always @(posedge H_count) begin
			in_cell = (H_count > H_SYNC + H_FRONT + H_SPAC + i*LIN_THCK + (i-1)* H_CELL_THCK &&
			H_count < H_SYNC + H_FRONT + H_SPAC + i*(LIN_THCK + H_CELL_THCK) &&
			V_count > V_SYNC + V_FRONT + V_TOP_SPAC + j*LIN_THCK + (j-1)* V_CELL_THCK &&
			V_count < V_SYNC + V_FRONT + V_TOP_SPAC + j*(LIN_THCK + V_CELL_THCK)) ? 1 : 0;
		
		H_dist = (H_count - H_SYNC - H_FRONT - H_SPAC - i*LIN_THCK - (i-1/2)*H_CELL_THCK + 22) * 
					(H_count - H_SYNC - H_FRONT - H_SPAC - i*LIN_THCK - (i-1/2)*H_CELL_THCK + 22);
		V_dist = (V_count - V_SYNC - V_FRONT - V_TOP_SPAC - j*LIN_THCK - (j-1/2)*V_CELL_THCK +15) * 
					(V_count - V_SYNC - V_FRONT - V_TOP_SPAC - j*LIN_THCK - (j-1/2)*V_CELL_THCK + 15);
		R_out <= in_cell && (H_dist + V_dist < 180) ? 8'b00000000 : 8'b00000000;
		G_out <= in_cell && (H_dist + V_dist < 180) ? 8'b00000000 : 8'b00000000;
		B_out <= in_cell && (H_dist + V_dist < 180) ? 8'b11111111 : 8'b00000000;
		
	end
	
endmodule



//---------------------FPGA Button Debounce Solution-------------------------

module debounce(clk, button_one, button_two, button_activity, button_one_out, button_two_out,button_activity_out);
input clk, button_one, button_two, button_activity;
reg [3:0] button_one_counter, button_two_counter, button_activity_counter;
output reg button_one_out, button_two_out, button_activity_out;
always @(posedge clk) begin
	if(~button_one && button_one_counter <3)begin // determining a threshold value which is 3
		button_one_counter <= button_one_counter +1;
		button_one_out <= 1;
		end
	else if(button_one) begin
		button_one_counter <= 0;
		button_one_out <=1;     //button one out is active low
		end
	else if(button_one_counter == 3)
		button_one_out = 0;
	
	
	if(~button_two && button_two_counter <3) begin
		button_two_counter <= button_two_counter +1;
		button_two_out <= 1;
		end
	if(button_two) begin
		button_two_counter <= 0;
		button_two_out <= 1;
		end
	if(button_two_counter == 3)
		button_two_out <= 0;
		
	if(~button_activity && button_activity_counter <3) begin
		button_activity_counter <= button_activity_counter +1;
		button_activity_out <= 1;
		end
	if(button_activity) begin
		button_activity_counter <= 0;
		button_activity_out <= 1;
		end
	if(button_activity_counter == 3)
		button_activity_out <= 0;
	end
endmodule




//-----------------------------Game Logic Part-------------------------

module controller(clk,button0_in,button1_in,act_in,H_Sync, V_Sync, divided_clk, R_out, G_out, B_out);

input clk,button0_in,button1_in,act_in;
output [7:0] R_out;
output [7:0] G_out;
output [7:0] B_out;
output wire divided_clk;
output wire H_Sync;
output wire V_Sync;

wire button0, button1, act;
reg [4:0] roundcount;
reg turn;
reg [3:0] drawcount;
reg [3:0] triwincount;
reg [3:0] circwincount;
reg error;
reg [299:0] arrayout;

reg [2:0] array[0:15][0:15];

reg [3:0] count;
reg [7:0] coordinate;
reg [7:0] recordval11;
reg [7:0] recordval12;
reg [7:0] recordval23;
reg [7:0] recordval24;
reg [7:0] cordwin;
reg [1:0] wld;
reg [2:0] insider;
reg cond;

integer i;
integer j;
integer k;
integer l;
integer m;
integer n;
integer insidecount;
reg [27:0] tcounter;

initial begin
	turn = 0;
	drawcount = 4'b0000;
	triwincount = 4'b0000;
	circwincount = 4'b0000;
	error = 0;
	count = 4'b0000;
	roundcount = 5'b00000;
	coordinate = 8'b00000000;
	wld = 2'b00;
	insidecount = 0;
	insider = 0;
	arrayout = 0;
	cond = 0;
	tcounter = 0;
	
	for (i=0;i<16;i=i+1) begin
		for (j=0;j<16;j=j+1) begin
			array[i][j] = 3'b000;
		end
	end
end

debounce(.clk(clk), .button_one(button0_in),.button_two(button1_in),
	.button_activity(act_in), .button_one_out(button0), .button_two_out(button1),
	.button_activity_out(act));

vga_display disp(.divided_clk(divided_clk), .V_Sync(V_Sync),
	.H_Sync(H_Sync), .board(arrayout), .R_out(R_out), .G_out(G_out),
	.B_out(B_out), .turn(turn), .wld(wld), .roundcount(roundcount), .triwincount(triwincount), 
	.circwincount(circwincount), .error(error));
	
clock_divider div (.clk(clk), .divided_clk(divided_clk));

always @(posedge divided_clk) begin
	if (count < 4'b1000) begin
		if (button0 == 0 && act == 1 && insidecount == 0) begin
			count <= count +1;
			insidecount <= 1;
			coordinate <= {1'b0,coordinate[7:1]};
		end
		else if (button1 ==0 && act ==1 && insidecount == 0) begin
			count <= count +1;
			coordinate <= {1'b1,coordinate[7:1]};
			insidecount <= 1;
		end
	end
	
	if ( button0 == 1 && button1 == 1 && act == 1) begin
		insidecount <= 0;
	end
	
	else if (count ==8 && act ==0 ) begin
		if (turn == 0 && array[coordinate[7:4] + 4'b0011][coordinate[3:0] + 4'b0011] == 3'b000 ) begin
			array[coordinate[7:4] + 4'b0011][coordinate[3:0] + 4'b0011] <= 3'b001;
			count <= 0;
			error <= 0;
			turn <= ~turn;
			cordwin <= {coordinate[3:0],coordinate[7:4]};
			roundcount <= roundcount +1;
			
			if ( roundcount == 5'b01010) begin
				array[recordval11[7:4]+ 4'b0011][recordval11[3:0]+4'b0011] <= 3'b011;
			end
			else if ( roundcount == 5'b01011) begin
				array[recordval12[7:4]+ 4'b0011][recordval12[3:0]+4'b0011] <= 3'b011;
			end
			else if ( roundcount == 5'b10110) begin
				array[recordval23[7:4]+ 4'b0011][recordval23[3:0]+4'b0011] <= 3'b011;
			end
			else if ( roundcount == 5'b10111) begin
				array[recordval24[7:4]+ 4'b0011][recordval24[3:0]+4'b0011] <= 3'b011;
			end
			
		end
		else if (turn ==1 && array[coordinate[7:4] + 4'b0011][coordinate[3:0] + 4'b0011] == 3'b000) begin
			array[coordinate[7:4] + 4'b0011][coordinate[3:0] + 4'b0011] <= 3'b010;
			count <= 0;
			error <= 0;
			turn <= ~turn;
			cordwin <= {coordinate[3:0],coordinate[7:4]};
			roundcount <= roundcount +1;
			
			if ( roundcount == 5'b01010) begin
				array[recordval11[7:4]+ 4'b0011][recordval11[3:0]+4'b0011] <= 3'b011;
			end
			else if ( roundcount == 5'b01011) begin
				array[recordval12[7:4]+ 4'b0011][recordval12[3:0]+4'b0011] <= 3'b011;
			end
			else if ( roundcount == 5'b10110) begin
				array[recordval23[7:4]+ 4'b0011][recordval23[3:0]+4'b0011] <= 3'b011;
			end
			else if ( roundcount == 5'b10111) begin
				array[recordval24[7:4]+ 4'b0011][recordval24[3:0]+4'b0011] <= 3'b011;
			end
		end
		else if ( array[coordinate[7:4] + 4'b0011][coordinate[3:0] + 4'b0011] != 3'b000) begin
			count <= 0;
			error <= 1;
		end
	end	
			
	if (roundcount == 5'b00001 && count ==0) begin
		recordval11 <= coordinate;
	end
	
	else if (roundcount == 5'b00010 && count ==0) begin
		recordval12 <= coordinate;
	end
	
	else if (roundcount == 5'b00011 && count ==0) begin
		recordval23 <= coordinate;
	end
	
	else if (roundcount == 5'b00100 && count ==0) begin
		recordval24 <= coordinate;
	end
	
	
	if (((array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0010][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0001][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0]][cordwin[7:4]+4'b0011] == 3'b001) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0010][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0001][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0100][cordwin[7:4]+4'b0011] == 3'b001) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0010][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0100][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0101][cordwin[7:4]+4'b0011] == 3'b001) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0100][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0101][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0110][cordwin[7:4]+4'b0011] == 3'b001) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0010] == 3'b001 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0001] == 3'b001 && array[cordwin[3:0] +4'b0011][cordwin[7:4]] == 3'b001) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0001] == 3'b001 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0010] == 3'b001 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0100] == 3'b001) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0010] == 3'b001 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0100] == 3'b001 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0101] == 3'b001) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0100] == 3'b001 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0101] == 3'b001 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0110] == 3'b001) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0010][cordwin[7:4]+4'b0010] == 3'b001 &&  array[cordwin[3:0] +4'b0001][cordwin[7:4]+4'b0001] == 3'b001 && array[cordwin[3:0]][cordwin[7:4]] == 3'b001) || ( array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0010][cordwin[7:4]+4'b0010] == 3'b001 && array[cordwin[3:0] +4'b0001][cordwin[7:4]+4'b0001] == 3'b001 && array[cordwin[3:0] +4'b0100][cordwin[7:4]+4'b0100] == 3'b001) || ( array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0010][cordwin[7:4]+4'b0010] == 3'b001 && array[cordwin[3:0] +4'b0100][cordwin[7:4]+4'b0100] == 3'b001 && array[cordwin[3:0] +4'b0101][cordwin[7:4]+4'b0101] == 3'b001) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0100][cordwin[7:4]+4'b0100] == 3'b001 && array[cordwin[3:0] +4'b0101][cordwin[7:4]+4'b0101] == 3'b001 && array[cordwin[3:0] +4'b0110][cordwin[7:4]+4'b0110] == 3'b001) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0010][cordwin[7:4]+4'b0100] == 3'b001 && array[cordwin[3:0] +4'b0001][cordwin[7:4]+4'b0101] == 3'b001 && array[cordwin[3:0]][cordwin[7:4]+4'b0110] == 3'b001) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0010][cordwin[7:4]+4'b0100] == 3'b001 && array[cordwin[3:0] +4'b0001][cordwin[7:4]+4'b0101] == 3'b001 && array[cordwin[3:0] +4'b0100][cordwin[7:4]+4'b0010] == 3'b001) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0010][cordwin[7:4]+4'b0100] == 3'b001 && array[cordwin[3:0] +4'b0100][cordwin[7:4]+4'b0010] == 3'b001 && array[cordwin[3:0] +4'b0101][cordwin[7:4]+4'b0001] == 3'b001) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b001 && array[cordwin[3:0] +4'b0100][cordwin[7:4]+4'b0010] == 3'b001 && array[cordwin[3:0] +4'b0101][cordwin[7:4]+4'b0001] == 3'b001 && array[cordwin[3:0] +4'b0110][cordwin[7:4]] == 3'b001)) && (cond == 0)) begin
		triwincount <= triwincount +1;
		wld <= 2'b01;
		cond <= 1;
	end
	else if (((array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0010][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0001][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0]][cordwin[7:4]+4'b0011] == 3'b010) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0010][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0001][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0100][cordwin[7:4]+4'b0011] == 3'b010) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0010][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0100][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0101][cordwin[7:4]+4'b0011] == 3'b010) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0100][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0101][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0110][cordwin[7:4]+4'b0011] == 3'b010) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0010] == 3'b010 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0001] == 3'b010 && array[cordwin[3:0] +4'b0011][cordwin[7:4]] == 3'b010) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0001] == 3'b010 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0010] == 3'b010 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0100] == 3'b010) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0010] == 3'b010 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0100] == 3'b010 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0101] == 3'b010) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0100] == 3'b010 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0101] == 3'b010 && array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0110] == 3'b010) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0010][cordwin[7:4]+4'b0010] == 3'b010 &&  array[cordwin[3:0] +4'b0001][cordwin[7:4]+4'b0001] == 3'b010 && array[cordwin[3:0]][cordwin[7:4]] == 3'b010) || ( array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0010][cordwin[7:4]+4'b0010] == 3'b010 && array[cordwin[3:0] +4'b0001][cordwin[7:4]+4'b0001] == 3'b010 && array[cordwin[3:0] +4'b0100][cordwin[7:4]+4'b0100] == 3'b010) || ( array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0010][cordwin[7:4]+4'b0010] == 3'b010 && array[cordwin[3:0] +4'b0100][cordwin[7:4]+4'b0100] == 3'b010 && array[cordwin[3:0] +4'b0101][cordwin[7:4]+4'b0101] == 3'b010) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0100][cordwin[7:4]+4'b0100] == 3'b010 && array[cordwin[3:0] +4'b0101][cordwin[7:4]+4'b0101] == 3'b010 && array[cordwin[3:0] +4'b0110][cordwin[7:4]+4'b0110] == 3'b010) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0010][cordwin[7:4]+4'b0100] == 3'b010 && array[cordwin[3:0] +4'b0001][cordwin[7:4]+4'b0101] == 3'b010 && array[cordwin[3:0]][cordwin[7:4]+4'b0110] == 3'b010) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0010][cordwin[7:4]+4'b0100] == 3'b010 && array[cordwin[3:0] +4'b0001][cordwin[7:4]+4'b0101] == 3'b010 && array[cordwin[3:0] +4'b0100][cordwin[7:4]+4'b0010] == 3'b010) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0010][cordwin[7:4]+4'b0100] == 3'b010 && array[cordwin[3:0] +4'b0100][cordwin[7:4]+4'b0010] == 3'b010 && array[cordwin[3:0] +4'b0101][cordwin[7:4]+4'b0001] == 3'b010) || (array[cordwin[3:0] +4'b0011][cordwin[7:4]+4'b0011] == 3'b010 && array[cordwin[3:0] +4'b0100][cordwin[7:4]+4'b0010] == 3'b010 && array[cordwin[3:0] +4'b0101][cordwin[7:4]+4'b0001] == 3'b010 && array[cordwin[3:0] +4'b0110][cordwin[7:4]] == 3'b010)) && (cond == 0)) begin
		circwincount <= circwincount +1;
		wld <= 2'b10;
		cond <= 1;
	end
	else if (roundcount == 25 && cond == 0) begin
		drawcount <= drawcount +1;
		wld <= 2'b11;
		cond <= 1;
		
	end
	
	if (cond == 1) begin
		tcounter <= tcounter +1;
		if (tcounter == 28'b1110111001101011001010000000 && (wld != 2'b11) ) begin
			tcounter <= 0;
			cond <= 0;
			wld <= 2'b00;
			roundcount <= 0;
			count <= 0;
			turn <= ~turn;
			for (k=0;k<16;k=k+1) begin
				for (l=0;l<16;l=l+1) begin
				array[l][k] = 3'b000;
				end
			end
		end
		else if (tcounter == 28'b1110111001101011001010000000 && (wld == 2'b11) ) begin
			tcounter <= 0;
			cond <= 0;
			wld <= 2'b00;
			roundcount <= 0;
			count <= 0;
			turn <= 0;
			for (k=0;k<16;k=k+1) begin
				for (l=0;l<16;l=l+1) begin
				array[l][k] = 3'b000;
				end
			end
		end
	end
		
end


always @* begin

	for (m=3;m<13;m=m+1) begin
		for (n=3;n<13;n=n+1) begin
			insider = {array[m][n][0],array[m][n][1],array[m][n][2]};
			arrayout = {insider,arrayout[299:3]};
		end
	end
end

endmodule
